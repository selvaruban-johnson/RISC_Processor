`include "risc_packet.sv"
`include "risc_generator.sv"
`include "risc_driver.sv"
`include "dut_if.sv"
`include "instruction_decodr.v"
`include "RISC.v"
`include "probe_packet.sv"
`include "probe_intf.sv"
//`include "risc_monitor.sv"
//`include "risc_alu_monitor.sv"
`include "risc_ram_monitor.sv"
`include "risc_coverage.sv"
//`include "risc_scoreboard.sv"
//`include "risc_alu_scoreboard.sv"
`include "risc_ram_scoreboard.sv"
`include "risc_environment.sv"
`include "risc_test.sv"
